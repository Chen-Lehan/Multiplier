`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2021/09/15 12:11:30
// Design Name: 
// Module Name: multiplier
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module multiplier(
    input   [31: 0]     X,
    input   [31: 0]     Y,
    output  [63: 0]     result
    );
    
    wire    [31: 0]     P_32    [15: 0];
    wire    [63: 0]     P_64    [15: 0];
    wire    [15: 0]     Cout_to_switch;
    wire    [15: 0]     Cout_to_wallacetree;
    wire    [15: 0]     N_64    [63: 0];
    wire    [63: 0]     src1;
    wire    [63: 0]     src2;
    wire    [63: 0]     C;
    wire    [63: 0]     S;
    wire                Cin;
    
    genvar i;
    generate
        for(i = 0; i < 32; i = i + 2) begin: booth_selector
            case(i)
                1: begin
                    booth_selector booth_selector(
                        .y0(             1'b0),
                        .y1(             Y[0]),
                        .y2(             Y[1]),
                        .X (                X),
                        .P (          P_32[0]),
                        .C (Cout_to_switch[0])
                    );
                end
                
                default: begin
                    booth_selector booth_selector(
                        .y0(           Y[i - 1]),
                        .y1(               Y[i]),
                        .y2(           Y[i + 1]),
                        .X (                  X),
                        .P (          P_32[i/2]),
                        .C (Cout_to_switch[i/2])
                    );
                end
             endcase
        end
    endgenerate
    
    assign P_64[0] = {{32{P_32[0][31]}},
                          P_32[0]
                     };
    assign P_64[1] = {{30{P_32[1][31]}},
                          P_32[1],
                      { 2{P_32[1][31]}}
                     };
    assign P_64[2] = {{28{P_32[2][31]}},
                          P_32[2],
                      { 4{P_32[2][31]}}
                     };
    assign P_64[3] = {{26{P_32[3][31]}},
                          P_32[3],
                      { 6{P_32[3][31]}}
                     };
    assign P_64[4] = {{24{P_32[4][31]}},
                          P_32[4],
                      { 8{P_32[4][31]}}
                     };
    assign P_64[5] = {{22{P_32[5][31]}},
                          P_32[5],
                      {10{P_32[5][31]}}
                     };
    assign P_64[6] = {{20{P_32[6][31]}},
                          P_32[6],
                      {12{P_32[6][31]}}
                     };
    assign P_64[7] = {{18{P_32[7][31]}},
                          P_32[7],
                      {14{P_32[7][31]}}
                     };
    assign P_64[8] = {{16{P_32[8][31]}},
                          P_32[8],
                      {16{P_32[8][31]}}
                     };
    assign P_64[9] = {{14{P_32[9][31]}},
                          P_32[9],
                      {18{P_32[9][31]}}
                     };
    assign P_64[10] = {{12{P_32[10][31]}},
                           P_32[10],
                       {20{P_32[10][31]}}
                     };
    assign P_64[11] = {{10{P_32[11][31]}},
                           P_32[11],
                       {22{P_32[11][31]}}
                     };
    assign P_64[12] = {{ 8{P_32[12][31]}},
                           P_32[12],
                       {24{P_32[12][31]}}
                     };
    assign P_64[13] = {{ 6{P_32[13][31]}},
                           P_32[13],
                       {26{P_32[13][31]}}
                     };
    assign P_64[14] = {{ 4{P_32[14][31]}},
                           P_32[14],
                       {28{P_32[14][31]}}
                     };
    assign P_64[15] = {{ 2{P_32[15][31]}},
                           P_32[15],
                       {30{P_32[15][31]}}
                     };
                     
    
    switch switch(
        .P_0(P_64[0]),
        .P_1(P_64[1]),
        .P_2(P_64[2]),
        .P_3(P_64[3]),
        .P_4(P_64[4]),
        .P_5(P_64[5]),
        .P_6(P_64[6]),
        .P_7(P_64[7]),
        .P_8(P_64[8]),
        .P_9(P_64[9]),
        .P_10(P_64[10]),
        .P_11(P_64[11]),
        .P_12(P_64[12]),
        .P_13(P_64[13]),
        .P_14(P_64[14]),
        .P_15(P_64[15]),
        .Cin(Cout_to_switch),
        .N_0(N_64[0]),
        .N_1(N_64[1]),
        .N_2(N_64[2]),
        .N_3(N_64[3]),
        .N_4(N_64[4]),
        .N_5(N_64[5]),
        .N_6(N_64[6]),
        .N_7(N_64[7]),
        .N_8(N_64[8]),
        .N_9(N_64[9]),
        .N_10(N_64[10]),
        .N_11(N_64[11]),
        .N_12(N_64[12]),
        .N_13(N_64[13]),
        .N_14(N_64[14]),
        .N_15(N_64[15]),
        .N_16(N_64[16]),
        .N_17(N_64[17]),
        .N_18(N_64[18]),
        .N_19(N_64[19]),
        .N_20(N_64[20]),
        .N_21(N_64[21]),
        .N_22(N_64[22]),
        .N_23(N_64[23]),
        .N_24(N_64[24]),
        .N_25(N_64[25]),
        .N_26(N_64[26]),
        .N_27(N_64[27]),
        .N_28(N_64[28]),
        .N_29(N_64[29]),
        .N_30(N_64[30]),
        .N_31(N_64[31]),
        .N_32(N_64[32]),
        .N_33(N_64[33]),
        .N_34(N_64[34]),
        .N_35(N_64[35]),
        .N_36(N_64[36]),
        .N_37(N_64[37]),
        .N_38(N_64[38]),
        .N_39(N_64[39]),
        .N_40(N_64[40]),
        .N_41(N_64[41]),
        .N_42(N_64[42]),
        .N_43(N_64[43]),
        .N_44(N_64[44]),
        .N_45(N_64[45]),
        .N_46(N_64[46]),
        .N_47(N_64[47]),
        .N_48(N_64[48]),
        .N_49(N_64[49]),
        .N_50(N_64[50]),
        .N_51(N_64[51]),
        .N_52(N_64[52]),
        .N_53(N_64[53]),
        .N_54(N_64[54]),
        .N_55(N_64[55]),
        .N_56(N_64[56]),
        .N_57(N_64[57]),
        .N_58(N_64[58]),
        .N_59(N_64[59]),
        .N_60(N_64[60]),
        .N_61(N_64[61]),
        .N_62(N_64[62]),
        .N_63(N_64[63]),
        .Cout(Cout_to_wallacetree)
    );
    
    wallace_tree wallace_tree(
        
        .N_0(N_64[0]),
        .N_1(N_64[1]),
        .N_2(N_64[2]),
        .N_3(N_64[3]),
        .N_4(N_64[4]),
        .N_5(N_64[5]),
        .N_6(N_64[6]),
        .N_7(N_64[7]),
        .N_8(N_64[8]),
        .N_9(N_64[9]),
        .N_10(N_64[10]),
        .N_11(N_64[11]),
        .N_12(N_64[12]),
        .N_13(N_64[13]),
        .N_14(N_64[14]),
        .N_15(N_64[15]),
        .N_16(N_64[16]),
        .N_17(N_64[17]),
        .N_18(N_64[18]),
        .N_19(N_64[19]),
        .N_20(N_64[20]),
        .N_21(N_64[21]),
        .N_22(N_64[22]),
        .N_23(N_64[23]),
        .N_24(N_64[24]),
        .N_25(N_64[25]),
        .N_26(N_64[26]),
        .N_27(N_64[27]),
        .N_28(N_64[28]),
        .N_29(N_64[29]),
        .N_30(N_64[30]),
        .N_31(N_64[31]),
        .N_32(N_64[32]),
        .N_33(N_64[33]),
        .N_34(N_64[34]),
        .N_35(N_64[35]),
        .N_36(N_64[36]),
        .N_37(N_64[37]),
        .N_38(N_64[38]),
        .N_39(N_64[39]),
        .N_40(N_64[40]),
        .N_41(N_64[41]),
        .N_42(N_64[42]),
        .N_43(N_64[43]),
        .N_44(N_64[44]),
        .N_45(N_64[45]),
        .N_46(N_64[46]),
        .N_47(N_64[47]),
        .N_48(N_64[48]),
        .N_49(N_64[49]),
        .N_50(N_64[50]),
        .N_51(N_64[51]),
        .N_52(N_64[52]),
        .N_53(N_64[53]),
        .N_54(N_64[54]),
        .N_55(N_64[55]),
        .N_56(N_64[56]),
        .N_57(N_64[57]),
        .N_58(N_64[58]),
        .N_59(N_64[59]),
        .N_60(N_64[60]),
        .N_61(N_64[61]),
        .N_62(N_64[62]),
        .N_63(N_64[63]),
        .Cin(Cout_to_wallacetree[13:0]),
        .C(C),
        .S(S)
    );
    
    assign src1 = {C[62:0], Cout_to_wallacetree[14]};
    assign src2 = S;
    assign Cin  = Cout_to_wallacetree[15];
    
    assign result = src1 + src2 + Cin;     
    
endmodule
